// PIEZO_BGMUSIC.sv

// C    16.35   32.70   65.41   130.81  261.63  523.25  1046.50 2093.00  4186.01
parameter C0 = 61162; // 16.35 Hz
parameter C1 = 30581; // 32.70 Hz
parameter C2 = 15288; // 65.41 Hz
parameter C3 = 7645; // 130.81 Hz
parameter C4 = 3822; // 261.63 Hz
parameter C5 = 1911; // 523.25 Hz
parameter C6 = 956; // 1046.50 Hz
parameter C7 = 478; // 2093.00 Hz
parameter C8 = 239; // 4186.01 Hz
// C#   17.32   34.65   69.30   138.59  277.18  554.37  1108.73 2217.46  4434.92
parameter C_s0 = 57737; // 17.32 Hz
parameter C_s1 = 28860; // 34.65 Hz
parameter C_s2 = 14430; // 69.30 Hz
parameter C_s3 = 7216; // 138.59 Hz
parameter C_s4 = 3608; // 277.18 Hz
parameter C_s5 = 1804; // 554.37 Hz
parameter C_s6 = 902; // 1108.73 Hz
parameter C_s7 = 451; // 2217.46 Hz
parameter C_s8 = 225; // 4434.92 Hz
// D    18.35   36.71   73.42   146.83  293.66  587.33  1174.66 2349.32  4698.64
parameter D0 = 54496; // 18.35 Hz
parameter D1 = 27241; // 36.71 Hz
parameter D2 = 13620; // 73.42 Hz
parameter D3 = 6811; // 146.83 Hz
parameter D4 = 3405; // 293.66 Hz
parameter D5 = 1703; // 587.33 Hz
parameter D6 = 851; // 1174.66 Hz
parameter D7 = 426; // 2349.32 Hz
parameter D8 = 213; // 4698.64 Hz
// D#   19.45   38.89   77.78   155.56  311.13  622.25  1244.51 2489.02  4978.03
parameter D_s0 = 51414; // 19.45 Hz
parameter D_s1 = 25714; // 38.89 Hz
parameter D_s2 = 12857; // 77.78 Hz
parameter D_s3 = 6428; // 155.56 Hz
parameter D_s4 = 3214; // 311.13 Hz
parameter D_s5 = 1607; // 622.25 Hz
parameter D_s6 = 804; // 1244.51 Hz
parameter D_s7 = 402; // 2489.02 Hz
parameter D_s8 = 201; // 4978.03 Hz
// E    20.60   41.20   82.41   164.81  329.63  659.26  1318.51 2637.02  5274.04
parameter E0 = 48544; // 20.60 Hz
parameter E1 = 24272; // 41.20 Hz
parameter E2 = 12134; // 82.41 Hz
parameter E3 = 6068; // 164.81 Hz
parameter E4 = 3034; // 329.63 Hz
parameter E5 = 1517; // 659.26 Hz
parameter E6 = 758; // 1318.51 Hz
parameter E7 = 379; // 2637.02 Hz
parameter E8 = 190; // 5274.04 Hz
// F    21.83   43.65   87.31   174.61  349.23  698.46  1396.91 2793.83  5587.65
parameter F0 = 45809; // 21.83 Hz
parameter F1 = 22910; // 43.65 Hz
parameter F2 = 11453; // 87.31 Hz
parameter F3 = 5727; // 174.61 Hz
parameter F4 = 2863; // 349.23 Hz
parameter F5 = 1432; // 698.46 Hz
parameter F6 = 716; // 1396.91 Hz
parameter F7 = 358; // 2793.83 Hz
parameter F8 = 179; // 5587.65 Hz
// F#   23.12   46.25   92.50   185.00  369.99  739.99  1479.98 2959.96  5919.91
parameter F_s0 = 43253; // 23.12 Hz
parameter F_s1 = 21622; // 46.25 Hz
parameter F_s2 = 10811; // 92.50 Hz
parameter F_s3 = 5405; // 185.00 Hz
parameter F_s4 = 2703; // 369.99 Hz
parameter F_s5 = 1351; // 739.99 Hz
parameter F_s6 = 676; // 1479.98 Hz
parameter F_s7 = 338; // 2959.96 Hz
parameter F_s8 = 169; // 5919.91 Hz
// G    24.50   49.00   98.00   196.00  392.00  783.99  1567.98 3135.96  6271.93
parameter G0 = 40816; // 24.50 Hz
parameter G1 = 20408; // 49.00 Hz
parameter G2 = 10204; // 98.00 Hz
parameter G3 = 5102; // 196.00 Hz
parameter G4 = 2551; // 392.00 Hz
parameter G5 = 1276; // 783.99 Hz
parameter G6 = 638; // 1567.98 Hz
parameter G7 = 319; // 3135.96 Hz
parameter G8 = 159; // 6271.93 Hz
// G#   25.96   51.91   103.83  207.65  415.30  830.61  1661.22 3322.44  6644.88
parameter G_s0 = 38521; // 25.96 Hz
parameter G_s1 = 19264; // 51.91 Hz
parameter G_s2 = 9631; // 103.83 Hz
parameter G_s3 = 4816; // 207.65 Hz
parameter G_s4 = 2408; // 415.30 Hz
parameter G_s5 = 1204; // 830.61 Hz
parameter G_s6 = 602; // 1661.22 Hz
parameter G_s7 = 301; // 3322.44 Hz
parameter G_s8 = 150; // 6644.88 Hz
// A    27.50   55.00   110.00  220.00  440.00  880.00  1760.00 3520.00  7040.00
parameter A0 = 36364; // 27.50 Hz
parameter A1 = 18182; // 55.00 Hz
parameter A2 = 9091; // 110.00 Hz
parameter A3 = 4545; // 220.00 Hz
parameter A4 = 2273; // 440.00 Hz
parameter A5 = 1136; // 880.00 Hz
parameter A6 = 568; // 1760.00 Hz
parameter A7 = 284; // 3520.00 Hz
parameter A8 = 142; // 7040.00 Hz
// A#   29.14   58.27   116.54  233.08  466.16  932.33  1864.66 3729.31  7458.62
parameter A_s0 = 34317; // 29.14 Hz
parameter A_s1 = 17161; // 58.27 Hz
parameter A_s2 = 8581; // 116.54 Hz
parameter A_s3 = 4290; // 233.08 Hz
parameter A_s4 = 2145; // 466.16 Hz
parameter A_s5 = 1073; // 932.33 Hz
parameter A_s6 = 536; // 1864.66 Hz
parameter A_s7 = 268; // 3729.31 Hz
parameter A_s8 = 134; // 7458.62 Hz
// B    30.87   61.74   123.47  246.94  493.88  987.77  1975.53 3951.07  7902.13
parameter B0 = 32394; // 30.87 Hz
parameter B1 = 16197; // 61.74 Hz
parameter B2 = 8099; // 123.47 Hz
parameter B3 = 4050; // 246.94 Hz
parameter B4 = 2025; // 493.88 Hz
parameter B5 = 1012; // 987.77 Hz
parameter B6 = 506; // 1975.53 Hz
parameter B7 = 253; // 3951.07 Hz
parameter B8 = 127; // 7902.13 Hz

parameter PAUSE = -10;
parameter ENDL = -1;

typedef struct {
    int tone;
    int sstart;
    int llast;
} note;

parameter length_of_ballgame = 239;
parameter length_of_dearX = 108;
parameter length_of_narco = 280;

parameter note ballgame[238:0] = {'{C4, 0, 242718}, '{PAUSE, 242719, 582523}, '{C5, 582524, 825242}, '{PAUSE, 825243, 873785}, '{A4, 873786, 1116504}, '{PAUSE, 1116505, 1165047}, '{G4, 1165048, 1407766}, '{PAUSE, 1407767, 1456309}, '{E4, 1456310, 1699028}, '{PAUSE, 1699029, 1747571}, '{G4, 1747572, 2548542}, '{PAUSE, 2548543, 2621357}, '{D4, 2621358, 3422328}, '{PAUSE, 3422329, 3495143}, '{C4, 3495144, 3737862}, '{PAUSE, 3737863, 4077667}, '{C5, 4077668, 4320386}, '{PAUSE, 4320387, 4368929}, '{A4, 4368930, 4611648}, '{PAUSE, 4611649, 4660191}, '{G4, 4660192, 4902910}, '{PAUSE, 4902911, 4951453}, '{E4, 4951454, 5194172}, '{PAUSE, 
5194173, 5242715}, '{G4, 5242716, 6626210}, '{PAUSE, 6626211, 6990287}, '{A4, 6990288, 7233006}, '{PAUSE, 7233007, 7281549}, '{G_s4, 7281550, 7524268}, '{PAUSE, 7524269, 7572811}, '{A4, 7572812, 7815530}, '{PAUSE, 7815531, 7864073}, '{E4, 7864074, 8106792}, '{PAUSE, 8106793, 8155335}, '{F4, 8155336, 8398054}, '{PAUSE, 8398055, 8446597}, '{G4, 8446598, 8689316}, '{PAUSE, 8689317, 8737859}, '{A4, 8737860, 8980578}, '{PAUSE, 8980579, 9320383}, '{F4, 9320384, 9563102}, '{PAUSE, 9563103, 9611645}, '{D4, 9611646, 10412616}, '{PAUSE, 10412617, 10485431}, '{A4, 10485432, 10728150}, '{PAUSE, 10728151, 11067955}, '{A4, 11067956, 11310674}, '{PAUSE, 11310675, 11359217}, '{A4, 11359218, 11601936}, '{PAUSE, 11601937, 11650479}, '{B4, 11650480, 11893198}, '{PAUSE, 11893199, 11941741}, '{C5, 11941742, 12184460}, '{PAUSE, 12184461, 12233003}, '{D5, 12233004, 12475722}, '{PAUSE, 12475723, 12524265}, '{B4, 12524266, 12766984}, '{PAUSE, 12766985, 12815527}, '{A4, 12815528, 13058246}, '{PAUSE, 13058247, 13106789}, '{G4, 13106790, 13349508}, '{PAUSE, 13349509, 13398051}, '{F4, 13398052, 13640770}, '{PAUSE, 13640771, 13689313}, '{D4, 13689314, 13932032}, '{PAUSE, 13932033, 13980575}, '{C4, 13980576, 14223294}, '{PAUSE, 14223295, 14563099}, '{C5, 14563100, 14805818}, '{PAUSE, 14805819, 14854361}, '{A4, 14854362, 15097080}, '{PAUSE, 15097081, 15145623}, '{G4, 15145624, 15388342}, '{PAUSE, 15388343, 15436885}, '{E4, 15436886, 15679604}, '{PAUSE, 15679605, 15728147}, '{G4, 15728148, 16529118}, '{PAUSE, 16529119, 16601933}, '{D4, 16601934, 17402904}, '{PAUSE, 17402905, 17475719}, '{C4, 17475720, 17718438}, '{PAUSE, 17718439, 18058243}, '{D4, 18058244, 18300962}, '{PAUSE, 18300963, 18349505}, '{E4, 18349506, 18592224}, '{PAUSE, 18592225, 18640767}, '{F4, 18640768, 18883486}, '{PAUSE, 18883487, 18932029}, '{G4, 18932030, 19174748}, '{PAUSE, 19174749, 19223291}, '{A4, 19223292, 20339796}, '{PAUSE, 20339797, 20388339}, '{A4, 20388340, 20631058}, '{PAUSE, 20631059, 20679601}, '{B4, 20679602, 20922320}, '{PAUSE, 20922321, 20970863}, '{C5, 20970864, 21213582}, '{PAUSE, 21213583, 21844649}, '{C5, 21844650, 22087368}, '{PAUSE, 22087369, 22718435}, '{C5, 22718436, 22961154}, '{PAUSE, 22961155, 23009697}, '{B4, 23009698, 23252416}, '{PAUSE, 23252417, 23300959}, '{A4, 23300960, 23543678}, '{PAUSE, 23543679, 23592221}, '{G4, 23592222, 23834940}, '{PAUSE, 23834941, 23883483}, '{F_s4, 23883484, 24126202}, '{PAUSE, 24126203, 24174745}, '{G4, 24174746, 24417464}, '{PAUSE, 24417465, 24466007}, '{A4, 24466008, 25266978}, '{PAUSE, 25266979, 25339793}, '{B4, 25339794, 26140764}, '{PAUSE, 26140765, 26213579}, '{C5, 26213580, 27888336}, '{PAUSE, 27888337, 27961151}, '{C4, 27961152, 28203870}, '{PAUSE, 28203871, 28543675}, '{C5, 28543676, 28786394}, '{PAUSE, 28786395, 28834937}, '{A4, 28834938, 29077656}, '{PAUSE, 29077657, 29126199}, '{G4, 29126200, 29368918}, '{PAUSE, 29368919, 29417461}, '{E4, 29417462, 29660180}, '{PAUSE, 29660181, 29708723}, '{G4, 29708724, 30509694}, '{PAUSE, 30509695, 30582509}, '{D4, 30582510, 31383480}, '{PAUSE, 31383481, 31456295}, '{C4, 31456296, 31699014}, '{PAUSE, 31699015, 32038819}, '{C5, 32038820, 32281538}, '{PAUSE, 32281539, 32330081}, '{A4, 32330082, 32572800}, '{PAUSE, 32572801, 32621343}, '{G4, 32621344, 32864062}, '{PAUSE, 32864063, 32912605}, '{E4, 32912606, 33155324}, '{PAUSE, 33155325, 33203867}, '{G4, 33203868, 34587362}, '{PAUSE, 34587363, 34660177}, '{G_s4, 34660178, 34902896}, '{PAUSE, 34902897, 34951439}, '{A4, 34951440, 35194158}, '{PAUSE, 35194159, 35242701}, '{G_s4, 35242702, 35485420}, '{PAUSE, 35485421, 35533963}, '{A4, 35533964, 35776682}, '{PAUSE, 35776683, 35825225}, '{E4, 35825226, 36067944}, '{PAUSE, 36067945, 36116487}, '{F4, 36116488, 36359206}, '{PAUSE, 36359207, 36407749}, '{G4, 36407750, 36650468}, '{PAUSE, 36650469, 36699011}, '{A4, 36699012, 36941730}, '{PAUSE, 36941731, 37281535}, '{F4, 37281536, 37524254}, '{PAUSE, 37524255, 37572797}, '{D4, 37572798, 38082506}, '{PAUSE, 38082507, 38446583}, '{A4, 38446584, 38956292}, '{PAUSE, 38956293, 39029107}, '{A4, 39029108, 39271826}, '{PAUSE, 39271827, 39320369}, '{A4, 39320370, 39563088}, '{PAUSE, 39563089, 39611631}, '{B4, 39611632, 39854350}, '{PAUSE, 39854351, 39902893}, '{C5, 39902894, 40145612}, '{PAUSE, 40145613, 40194155}, '{D5, 40194156, 40436874}, '{PAUSE, 40436875, 40485417}, '{B4, 40485418, 40728136}, '{PAUSE, 40728137, 40776679}, '{A4, 40776680, 41019398}, '{PAUSE, 41019399, 41067941}, '{G4, 41067942, 41310660}, '{PAUSE, 41310661, 41359203}, '{F4, 41359204, 41601922}, '{PAUSE, 41601923, 41650465}, '{D4, 41650466, 41893184}, '{PAUSE, 41893185, 41941727}, '{C4, 41941728, 
42184446}, '{PAUSE, 42184447, 42524251}, '{C5, 42524252, 42766970}, '{PAUSE, 42766971, 42815513}, '{A4, 42815514, 43058232}, '{PAUSE, 43058233, 43106775}, '{G4, 43106776, 43349494}, '{PAUSE, 43349495, 
43398037}, '{E4, 43398038, 43640756}, '{PAUSE, 43640757, 43689299}, '{G4, 43689300, 44490270}, '{PAUSE, 44490271, 44563085}, '{D4, 44563086, 45364056}, '{PAUSE, 45364057, 45436871}, '{C4, 45436872, 45946580}, '{PAUSE, 45946581, 46019395}, '{D4, 46019396, 46262114}, '{PAUSE, 46262115, 46310657}, '{E4, 46310658, 46553376}, '{PAUSE, 46553377, 46601919}, '{F4, 46601920, 46844638}, '{PAUSE, 46844639, 46893181}, '{G4, 46893182, 47135900}, '{PAUSE, 47135901, 47184443}, '{A4, 47184444, 48300948}, '{PAUSE, 48300949, 48349491}, '{A4, 48349492, 48592210}, '{PAUSE, 48592211, 48640753}, '{B4, 48640754, 48883472}, '{PAUSE, 48883473, 48932015}, '{C5, 48932016, 49174734}, '{PAUSE, 49174735, 49805801}, '{C5, 49805802, 50048520}, '{PAUSE, 50048521, 50679587}, '{C5, 50679588, 50922306}, '{PAUSE, 50922307, 50970849}, '{B4, 50970850, 51213568}, '{PAUSE, 51213569, 51262111}, '{A4, 51262112, 51504830}, '{PAUSE, 51504831, 51553373}, '{G4, 51553374, 51796092}, '{PAUSE, 51796093, 51844635}, '{F_s4, 51844636, 52087354}, '{PAUSE, 52087355, 52135897}, '{G4, 52135898, 52378616}, '{PAUSE, 52378617, 52427159}, '{A4, 52427160, 53228130}, '{PAUSE, 53228131, 53300945}, '{B4, 53300946, 54101916}, '{PAUSE, 54101917, 54174731}, '{C5, 54174732, 55291236}, '{PAUSE, 55291237, 57291237}, '{ENDL, 57291238, 57291248}};


parameter note dearX[107:0] = {'{A5, 0, 312500}, '{PAUSE, 312501, 319148}, '{G5, 319149, 631648}, '{PAUSE, 631649, 638296}, '{F_s5, 638297, 950797}, '{PAUSE, 950798, 957444}, '{A5, 957445, 1110371}, '{PAUSE, 1110372, 1117019}, '{A5, 1117020, 1429519}, '{PAUSE, 1429520, 1436167}, '{F_s5, 1436168, 1589094}, '{PAUSE, 1589095, 1595741}, '{F_s5, 1595742, 1908242}, '{PAUSE, 1908243, 1914890}, '{E5, 1914891, 2446805}, '{PAUSE, 2446806, 2553187}, '{A5, 2553188, 3085102}, '{PAUSE, 3085103, 3191484}, '{D6, 3191485, 3503985}, '{PAUSE, 3503986, 3510632}, '{C_s6, 3510633, 3663559}, '{PAUSE, 3663560, 3670207}, '{B5, 3670208, 4142282}, '{PAUSE, 4142283, 4148930}, '{A5, 4148931, 4301856}, '{PAUSE, 4301857, 4308504}, '{F_s5, 4308505, 4461430}, '{PAUSE, 4461431, 4468078}, '{F_s5, 4468079, 4999993}, '{PAUSE, 4999994, 5744672}, '{D5, 5744673, 6216747}, '{PAUSE, 6216748, 6223395}, '{E5, 6223396, 6695470}, '{PAUSE, 
6695471, 6702118}, '{F_s5, 6702119, 7014618}, '{PAUSE, 7014619, 7021266}, '{E5, 7021267, 7333767}, '{PAUSE, 7333768, 7340414}, '{D5, 7340415, 7493341}, '{PAUSE, 7493342, 7499989}, '{D5, 7499990, 8191478}, '{PAUSE, 8191479, 8297860}, '{G5, 8297861, 8610361}, '{PAUSE, 8610362, 8617008}, '{F_s5, 8617009, 8929509}, '{PAUSE, 8929510, 8936157}, '{G5, 8936158, 9089083}, '{PAUSE, 9089084, 9095731}, '{A5, 9095732, 9408232}, '{PAUSE, 9408233, 9414880}, '{E5, 9414881, 10106369}, '{PAUSE, 10106370, 10212751}, '{A5, 10212752, 10525252}, '{PAUSE, 10525253, 10531900}, '{G5, 10531901, 10844400}, '{PAUSE, 10844401, 10851048}, '{F_s5, 10851049, 11163549}, '{PAUSE, 11163550, 11170196}, '{A5, 11170197, 11323123}, '{PAUSE, 11323124, 11329771}, '{A5, 11329772, 11642271}, '{PAUSE, 11642272, 11648919}, '{F_s5, 11648920, 11801846}, '{PAUSE, 11801847, 11808493}, '{F_s5, 11808494, 12120994}, '{PAUSE, 12120995, 12127642}, '{E5, 12127643, 12659557}, '{PAUSE, 12659558, 12765939}, '{A5, 12765940, 13297854}, '{PAUSE, 13297855, 13404236}, 
'{D6, 13404237, 13716737}, '{PAUSE, 13716738, 13723384}, '{C_s6, 13723385, 13876311}, '{PAUSE, 13876312, 13882959}, '{B5, 13882960, 14355034}, '{PAUSE, 14355035, 14361682}, '{D6, 14361683, 14514608}, '{PAUSE, 14514609, 14521256}, '{A5, 14521257, 14674182}, '{PAUSE, 14674183, 14680830}, '{A5, 14680831, 15212745}, '{PAUSE, 15212746, 15957424}, '{D5, 15957425, 16429499}, '{PAUSE, 16429500, 16436147}, '{E5, 16436148, 16908222}, '{PAUSE, 16908223, 16914870}, '{F_s5, 16914871, 17227370}, '{PAUSE, 17227371, 17234018}, '{E5, 17234019, 17546519}, '{PAUSE, 17546520, 17553166}, '{D5, 17553167, 17706093}, '{PAUSE, 17706094, 17712741}, '{D5, 17712742, 18404230}, '{PAUSE, 18404231, 18510612}, '{G5, 18510613, 18663538}, '{PAUSE, 18663539, 18670186}, '{F_s5, 18670187, 18823113}, '{PAUSE, 18823114, 18829760}, '{E5, 18829761, 18982687}, '{PAUSE, 18982688, 18989335}, '{D5, 18989336, 19142261}, '{PAUSE, 19142262, 19148909}, '{E5, 19148910, 19461410}, '{PAUSE, 19461411, 19468057}, '{F_s5, 19468058, 19620984}, '{PAUSE, 19620985, 19627632}, '{D5, 19627633, 20319121}, '{PAUSE, 20319122, 22319121}};

parameter note narco[279:0] = {'{A5, 0, 400000}, '{PAUSE, 400001, 479999}, '{C5, 480000, 715000}, '{C6, 480000, 715000}, '{PAUSE, 715001, 719999}, '{D5, 720000, 955000}, '{D6, 720000, 955000}, '{PAUSE, 955001, 959999}, '{E5, 960000, 1360000}, '{E6, 960000, 1360000}, '{PAUSE, 1360001, 1919999}, '{E5, 1920000, 2275000}, '{E6, 1920000, 2275000}, '{PAUSE, 2275001, 2279999}, '{E5, 2280000, 2395000}, '{E6, 2280000, 2395000}, '{PAUSE, 2395001, 2399999}, '{D5, 2400000, 2635000}, '{D6, 2400000, 2635000}, '{PAUSE, 2635001, 2639999}, '{F5, 2640000, 2875000}, '{F6, 2640000, 2875000}, '{PAUSE, 2875001, 2879999}, '{E5, 2880000, 3280000}, '{E6, 2880000, 3280000}, '{PAUSE, 3280001, 3839999}, '{E5, 3840000, 4195000}, '{E6, 3840000, 4195000}, '{PAUSE, 4195001, 4199999}, '{E5, 4200000, 4315000}, '{E6, 4200000, 4315000}, '{PAUSE, 4315001, 4319999}, '{D5, 4320000, 4555000}, '{D6, 4320000, 4555000}, '{PAUSE, 4555001, 4559999}, '{F5, 4560000, 4795000}, '{F6, 4560000, 4795000}, '{PAUSE, 4795001, 4799999}, '{E5, 4800000, 5155000}, '{E6, 4800000, 5155000}, '{PAUSE, 5155001, 5159999}, '{E5, 5160000, 5275000}, '{E6, 5160000, 5275000}, '{PAUSE, 5275001, 5279999}, '{C5, 5280000, 5515000}, '{C6, 5280000, 5515000}, '{PAUSE, 5515001, 5519999}, '{B4, 5520000, 5755000}, '{B5, 5520000, 5755000}, '{PAUSE, 5755001, 5759999}, '{D5, 5760000, 6115000}, '{D6, 5760000, 6115000}, '{PAUSE, 6115001, 6119999}, '{D5, 6120000, 6235000}, '{D6, 6120000, 6235000}, '{PAUSE, 6235001, 6239999}, '{C5, 6240000, 6475000}, '{C6, 6240000, 6475000}, '{PAUSE, 6475001, 6479999}, '{B4, 6480000, 6715000}, '{B5, 6480000, 6715000}, '{PAUSE, 6715001, 6719999}, '{A4, 6720000, 7120000}, '{A5, 6720000, 7120000}, '{PAUSE, 7120001, 7679999}, '{A4, 7680000, 8080000}, '{A5, 7680000, 8080000}, '{PAUSE, 8080001, 8159999}, '{C5, 
8160000, 8395000}, '{C6, 8160000, 8395000}, '{PAUSE, 8395001, 8399999}, '{D5, 8400000, 8635000}, '{D6, 8400000, 8635000}, '{PAUSE, 8635001, 8639999}, '{E5, 8640000, 9040000}, '{E6, 8640000, 9040000}, '{PAUSE, 9040001, 9119999}, '{E5, 9120000, 9355000}, '{E6, 9120000, 9355000}, '{PAUSE, 9355001, 9359999}, '{E5, 9360000, 9595000}, '{E6, 9360000, 9595000}, '{PAUSE, 9595001, 9599999}, '{A5, 9600000, 9955000}, '{A6, 9600000, 9955000}, '{PAUSE, 9955001, 9959999}, '{A5, 9960000, 10075000}, '{A6, 9960000, 10075000}, '{PAUSE, 10075001, 10079999}, '{G5, 10080000, 10315000}, '{G6, 10080000, 10315000}, '{PAUSE, 10315001, 10319999}, '{F5, 10320000, 10555000}, '{F6, 10320000, 10555000}, '{PAUSE, 10555001, 10559999}, '{E5, 10560000, 10960000}, '{E6, 10560000, 10960000}, '{PAUSE, 10960001, 11279999}, '{E5, 11280000, 11515000}, '{E6, 11280000, 11515000}, '{PAUSE, 11515001, 11519999}, '{A5, 11520000, 11875000}, '{A6, 11520000, 11875000}, '{PAUSE, 11875001, 11879999}, '{A5, 11880000, 11995000}, '{A6, 11880000, 11995000}, '{PAUSE, 11995001, 11999999}, '{G5, 12000000, 12235000}, '{G6, 12000000, 12235000}, '{PAUSE, 12235001, 12239999}, '{F5, 12240000, 12475000}, '{F6, 12240000, 12475000}, '{PAUSE, 12475001, 12479999}, '{E5, 12480000, 12835000}, '{E6, 12480000, 12835000}, '{PAUSE, 12835001, 12839999}, '{E5, 12840000, 12955000}, '{E6, 12840000, 12955000}, '{PAUSE, 12955001, 12959999}, '{D5, 12960000, 13195000}, '{D6, 12960000, 13195000}, '{PAUSE, 13195001, 13199999}, '{C5, 13200000, 13435000}, '{C6, 13200000, 13435000}, '{PAUSE, 13435001, 13439999}, '{D5, 13440000, 13795000}, '{D6, 13440000, 13795000}, 
'{PAUSE, 13795001, 13799999}, '{D5, 13800000, 13915000}, '{D6, 13800000, 13915000}, '{PAUSE, 13915001, 13919999}, '{C5, 13920000, 14155000}, '{C6, 13920000, 14155000}, '{PAUSE, 14155001, 14159999}, '{B4, 14160000, 14395000}, '{B5, 14160000, 14395000}, '{PAUSE, 14395001, 14399999}, '{A4, 14400000, 14800000}, '{A5, 14400000, 14800000}, '{PAUSE, 14800001, 15359999}, '{A4, 15360000, 15760000}, '{A5, 15360000, 15760000}, '{PAUSE, 15760001, 15839999}, '{C5, 15840000, 16075000}, '{C6, 15840000, 16075000}, '{PAUSE, 16075001, 16079999}, '{D5, 16080000, 16315000}, '{D6, 16080000, 16315000}, '{PAUSE, 16315001, 16319999}, '{E5, 16320000, 16720000}, '{E6, 16320000, 16720000}, '{PAUSE, 16720001, 17279999}, '{E5, 17280000, 17635000}, '{E6, 17280000, 17635000}, '{PAUSE, 17635001, 17639999}, '{E5, 17640000, 17755000}, '{E6, 17640000, 17755000}, '{PAUSE, 17755001, 17759999}, '{D5, 
17760000, 17995000}, '{D6, 17760000, 17995000}, '{PAUSE, 17995001, 17999999}, '{F5, 18000000, 18235000}, '{F6, 18000000, 18235000}, '{PAUSE, 18235001, 18239999}, '{E5, 18240000, 18640000}, '{E6, 18240000, 18640000}, '{PAUSE, 18640001, 19199999}, '{E5, 19200000, 19555000}, '{E6, 19200000, 19555000}, '{PAUSE, 19555001, 19559999}, '{E5, 19560000, 19675000}, '{E6, 19560000, 19675000}, '{PAUSE, 19675001, 19679999}, '{D5, 19680000, 19915000}, '{D6, 19680000, 19915000}, '{PAUSE, 19915001, 19919999}, '{F5, 19920000, 20155000}, '{F6, 19920000, 20155000}, '{PAUSE, 20155001, 20159999}, '{E5, 20160000, 20515000}, '{E6, 20160000, 20515000}, '{PAUSE, 20515001, 20519999}, '{E5, 20520000, 20635000}, '{E6, 20520000, 20635000}, '{PAUSE, 20635001, 20639999}, '{C5, 20640000, 20875000}, '{C6, 20640000, 20875000}, '{PAUSE, 20875001, 20879999}, '{B4, 20880000, 21115000}, '{B5, 20880000, 21115000}, '{PAUSE, 21115001, 21119999}, '{D5, 21120000, 21475000}, '{D6, 21120000, 21475000}, '{PAUSE, 21475001, 21479999}, '{D5, 21480000, 21595000}, '{D6, 21480000, 21595000}, '{PAUSE, 21595001, 21599999}, '{C5, 21600000, 21835000}, '{C6, 21600000, 21835000}, '{PAUSE, 21835001, 21839999}, '{B4, 21840000, 22075000}, '{B5, 21840000, 22075000}, '{PAUSE, 22075001, 22079999}, '{A4, 22080000, 22480000}, '{A5, 22080000, 22480000}, '{PAUSE, 22480001, 23039999}, '{A4, 23040000, 23440000}, '{A5, 23040000, 23440000}, '{PAUSE, 23440001, 23519999}, '{C5, 23520000, 23755000}, '{C6, 23520000, 23755000}, '{PAUSE, 23755001, 23759999}, '{D5, 23760000, 23995000}, '{D6, 23760000, 23995000}, '{PAUSE, 23995001, 23999999}, '{E5, 24000000, 
24400000}, '{E6, 24000000, 24400000}, '{PAUSE, 24400001, 24479999}, '{E5, 24480000, 24715000}, '{E6, 24480000, 24715000}, '{PAUSE, 24715001, 24719999}, '{E5, 24720000, 24955000}, '{E6, 24720000, 24955000}, '{PAUSE, 24955001, 24959999}, '{A5, 24960000, 25315000}, '{A6, 24960000, 25315000}, '{PAUSE, 25315001, 25319999}, '{A5, 25320000, 25435000}, '{A6, 25320000, 25435000}, '{PAUSE, 25435001, 25439999}, '{G5, 25440000, 25675000}, '{G6, 25440000, 25675000}, '{PAUSE, 25675001, 25679999}, '{F5, 25680000, 25915000}, '{F6, 25680000, 25915000}, '{PAUSE, 25915001, 25919999}, '{E5, 25920000, 26320000}, '{E6, 25920000, 26320000}, '{PAUSE, 26320001, 26639999}, '{E5, 26640000, 26875000}, '{E6, 26640000, 26875000}, '{PAUSE, 26875001, 26879999}, '{A5, 26880000, 27235000}, '{A6, 26880000, 27235000}, '{PAUSE, 27235001, 27239999}, '{A5, 27240000, 27355000}, '{A6, 27240000, 27355000}, '{PAUSE, 27355001, 27359999}, '{G5, 27360000, 27595000}, '{G6, 27360000, 27595000}, '{PAUSE, 27595001, 27599999}, '{F5, 27600000, 27835000}, '{F6, 27600000, 27835000}, '{PAUSE, 27835001, 27839999}, '{E5, 27840000, 28195000}, '{E6, 27840000, 28195000}, '{PAUSE, 28195001, 28199999}, '{E5, 28200000, 28315000}, '{E6, 28200000, 28315000}, '{PAUSE, 28315001, 28319999}, '{D5, 28320000, 28555000}, '{D6, 28320000, 28555000}, '{PAUSE, 28555001, 28559999}, '{C5, 28560000, 28795000}, '{C6, 28560000, 28795000}, '{PAUSE, 28795001, 28799999}, '{D5, 28800000, 29155000}, '{D6, 28800000, 29155000}, '{PAUSE, 29155001, 29159999}, '{D5, 29160000, 29275000}, '{D6, 29160000, 29275000}, '{PAUSE, 29275001, 29279999}, '{C5, 29280000, 29515000}, '{C6, 29280000, 29515000}, '{PAUSE, 29515001, 29519999}, '{B4, 29520000, 29755000}, '{B5, 29520000, 29755000}, '{PAUSE, 29755001, 29759999}, '{A5, 29760000, 30160000}, '{PAUSE, 29760001, 31760001}};


parameter note christmas[743:0] = {'{G6, 0, 333333}, '{PAUSE, 333334, 399999}, '{B6, 400000, 845833}, '{PAUSE, 845834, 849999}, '{D7, 850000, 1245833}, '{PAUSE, 1245834, 1249999}, '{F_s7, 1250000, 1645833}, '{PAUSE, 1645834, 1649999}, '{G7, 1650000, 2045833}, '{PAUSE, 2045834, 2049999}, '{F_s7, 2050000, 2445833}, '{PAUSE, 2445834, 2449999}, '{D7, 2450000, 2795833}, '{PAUSE, 2795834, 2799999}, '{B6, 2800000, 3133333}, '{PAUSE, 3133334, 3199999}, '{G6, 3200000, 3533333}, '{PAUSE, 3533334, 3599999}, '{C7, 3600000, 3933333}, '{PAUSE, 3933334, 3999999}, '{D7, 4000000, 4445833}, '{PAUSE, 4445834, 4449999}, '{G7, 4450000, 4845833}, '{PAUSE, 4845834, 4849999}, '{D7, 4850000, 6300000}, '{PAUSE, 6300001, 6449999}, '{G4, 6450000, 8045833}, '{PAUSE, 8045834, 8049999}, '{B4, 8050000, 8545833}, '{PAUSE, 8545834, 8549999}, '{D5, 8550000, 9045833}, '{PAUSE, 9045834, 9049999}, '{F_s5, 9050000, 9545833}, '{PAUSE, 9545834, 9549999}, '{G5, 9550000, 9945833}, '{PAUSE, 9945834, 9949999}, '{F_s5, 9950000, 10445833}, '{PAUSE, 10445834, 10449999}, '{D5, 10450000, 11095833}, '{PAUSE, 11095834, 11099999}, '{E5, 11100000, 11495833}, '{PAUSE, 11495834, 11499999}, '{D5, 11500000, 12700000}, '{PAUSE, 12700001, 12849999}, '{A5, 12850000, 13395833}, '{PAUSE, 13395834, 13399999}, '{G5, 13400000, 13845833}, '{PAUSE, 13845834, 13849999}, '{F_s5, 13850000, 14145833}, '{PAUSE, 14145834, 14149999}, '{G5, 14150000, 14495833}, '{PAUSE, 14495834, 14499999}, '{F_s5, 14500000, 14895833}, '{PAUSE, 14895834, 14899999}, '{D5, 14900000, 15295833}, '{PAUSE, 15295834, 15299999}, '{E5, 15300000, 15695833}, '{PAUSE, 15695834, 15699999}, '{D5, 15700000, 16333333}, '{PAUSE, 16333334, 16749999}, '{C5, 16750000, 17095833}, '{PAUSE, 17095834, 17099999}, '{E5, 17100000, 17445833}, '{PAUSE, 17445834, 17449999}, '{G5, 17450000, 17895833}, '{PAUSE, 17895834, 17899999}, '{A5, 17900000, 18245833}, '{PAUSE, 18245834, 18249999}, '{B5, 18250000, 18645833}, '{PAUSE, 18645834, 18649999}, '{A5, 18650000, 19045833}, '{PAUSE, 19045834, 19049999}, '{G5, 19050000, 19395833}, '{PAUSE, 19395834, 19399999}, '{E5, 19400000, 19933333}, '{PAUSE, 19933334, 20349999}, '{B5, 20350000, 20695833}, '{PAUSE, 20695834, 20699999}, '{D6, 20700000, 20995833}, '{PAUSE, 20995834, 20999999}, '{B5, 21000000, 21533333}, '{PAUSE, 21533334, 21599999}, '{A5, 21600000, 21845833}, '{PAUSE, 21845834, 21849999}, '{B5, 21850000, 22145833}, '{PAUSE, 22145834, 22149999}, '{A5, 22150000, 22545833}, '{PAUSE, 22545834, 22549999}, '{G5, 22550000, 22995833}, '{PAUSE, 22995834, 22999999}, '{D_s5, 23000000, 23533333}, '{PAUSE, 23533334, 23949999}, '{G5, 23950000, 24295833}, '{PAUSE, 24295834, 24299999}, '{A5, 24300000, 24595833}, '{PAUSE, 24595834, 24599999}, '{F_s5, 24600000, 24945833}, '{PAUSE, 24945834, 24949999}, '{G5, 24950000, 25345833}, '{PAUSE, 25345834, 25349999}, '{E5, 25350000, 25745833}, '{PAUSE, 25745834, 25749999}, '{F_s5, 25750000, 26245833}, '{PAUSE, 26245834, 26249999}, '{D_s5, 26250000, 27533333}, '{PAUSE, 27533334, 28299999}, '{B5, 28300000, 28595833}, '{PAUSE, 28595834, 28599999}, '{A5, 28600000, 28945833}, '{PAUSE, 28945834, 28949999}, '{A5, 28950000, 29645833}, '{PAUSE, 29645834, 29649999}, '{G5, 29650000, 29945833}, '{PAUSE, 29945834, 29949999}, '{G5, 29950000, 30345833}, '{PAUSE, 30345834, 30349999}, '{A5, 30350000, 30745833}, '{PAUSE, 30745834, 30749999}, '{G5, 30750000, 31900000}, '{PAUSE, 31900001, 32799999}, '{D5, 32800000, 33145833}, '{PAUSE, 33145834, 33149999}, '{E5, 33150000, 33545833}, '{PAUSE, 33545834, 33549999}, '{G5, 33550000, 33945833}, '{PAUSE, 33945834, 33949999}, '{D6, 33950000, 34533333}, '{PAUSE, 34533334, 34599999}, '{C6, 34600000, 37133333}, '{PAUSE, 37133334, 38199999}, '{B5, 38200000, 39145833}, '{PAUSE, 39145834, 39149999}, '{A5, 39150000, 39895833}, '{PAUSE, 39895834, 39899999}, '{G5, 39900000, 40700000}, '{PAUSE, 40700001, 40799999}, '{E5, 40800000, 41445833}, '{PAUSE, 41445834, 41449999}, '{D_s5, 41450000, 42495833}, '{PAUSE, 42495834, 42499999}, '{A5, 42500000, 44300000}, '{PAUSE, 44300001, 44549999}, '{B5, 44550000, 46545833}, '{PAUSE, 46545834, 46549999}, '{A5, 46550000, 47445833}, '{PAUSE, 47445834, 47449999}, '{G5, 47450000, 51100000}, '{PAUSE, 51100001, 55999999}, '{G4, 56000000, 56333333}, '{PAUSE, 56333334, 56399999}, '{B4, 56400000, 56733333}, '{PAUSE, 56733334, 56799999}, '{D5, 56800000, 57133333}, '{PAUSE, 57133334, 57199999}, '{F_s5, 57200000, 57495833}, '{PAUSE, 57495834, 57499999}, '{G5, 57500000, 57895833}, '{PAUSE, 57895834, 57899999}, '{F_s5, 57900000, 58295833}, '{PAUSE, 58295834, 58299999}, '{E5, 58300000, 58695833}, 
'{PAUSE, 58695834, 58699999}, '{D5, 58700000, 59133333}, '{PAUSE, 59133334, 59199999}, '{A5, 59200000, 59533333}, '{PAUSE, 59533334, 59599999}, '{G5, 59600000, 59933333}, '{PAUSE, 59933334, 59999999}, '{G5, 60000000, 60333333}, '{PAUSE, 60333334, 60399999}, '{F_s5, 60400000, 60695833}, '{PAUSE, 60695834, 60699999}, '{G5, 60700000, 61095833}, '{PAUSE, 61095834, 61099999}, '{F_s5, 61100000, 61495833}, '{PAUSE, 61495834, 61499999}, '{E5, 61500000, 61895833}, '{PAUSE, 61895834, 61899999}, '{D5, 61900000, 62333333}, '{PAUSE, 62333334, 62399999}, '{C5, 62400000, 62733333}, '{PAUSE, 62733334, 62799999}, '{E5, 62800000, 63133333}, '{PAUSE, 63133334, 63199999}, '{G5, 63200000, 63533333}, '{PAUSE, 63533334, 63599999}, '{A5, 63600000, 63933333}, '{PAUSE, 63933334, 63999999}, '{B5, 64000000, 64333333}, '{PAUSE, 64333334, 64399999}, '{A5, 64400000, 64695833}, '{PAUSE, 64695834, 64699999}, '{G5, 64700000, 65095833}, '{PAUSE, 65095834, 65099999}, '{E5, 65100000, 65533333}, '{PAUSE, 65533334, 65599999}, '{C5, 65600000, 65933333}, '{PAUSE, 65933334, 65999999}, '{D_s5, 66000000, 66333333}, '{PAUSE, 66333334, 66399999}, '{G5, 66400000, 66733333}, '{PAUSE, 66733334, 66799999}, '{A5, 66800000, 67133333}, '{PAUSE, 67133334, 67199999}, '{A_s5, 67200000, 67533333}, '{PAUSE, 67533334, 67599999}, '{A5, 67600000, 67895833}, '{PAUSE, 67895834, 67899999}, '{G5, 67900000, 68700000}, '{PAUSE, 68700001, 68799999}, '{A5, 68800000, 69133333}, '{PAUSE, 69133334, 69199999}, '{G5, 69200000, 69495833}, '{PAUSE, 69495834, 69499999}, '{G5, 69500000, 69933333}, '{PAUSE, 69933334, 69999999}, '{F_s5, 70000000, 70295833}, 
'{PAUSE, 70295834, 70299999}, '{G5, 70300000, 70695833}, '{PAUSE, 70695834, 70699999}, '{F_s5, 70700000, 71095833}, '{PAUSE, 71095834, 71099999}, 
'{E5, 71100000, 71495833}, '{PAUSE, 71495834, 71499999}, '{D5, 71500000, 71933333}, '{PAUSE, 71933334, 71999999}, '{G4, 72000000, 72333333}, '{PAUSE, 72333334, 72399999}, '{B4, 72400000, 72733333}, '{PAUSE, 72733334, 72799999}, '{D5, 72800000, 73133333}, '{PAUSE, 73133334, 73199999}, '{F_s5, 73200000, 73495833}, '{PAUSE, 73495834, 73499999}, '{G5, 73500000, 73895833}, '{PAUSE, 73895834, 73899999}, '{F_s5, 73900000, 74295833}, '{PAUSE, 74295834, 74299999}, '{E5, 74300000, 75100000}, '{PAUSE, 75100001, 75599999}, '{B5, 75600000, 75895833}, '{PAUSE, 75895834, 75899999}, '{A5, 75900000, 75995833}, '{PAUSE, 75995834, 75999999}, '{B5, 76000000, 76333333}, '{PAUSE, 76333334, 76399999}, '{A5, 76400000, 76733333}, '{PAUSE, 76733334, 76799999}, '{B5, 76800000, 77133333}, '{PAUSE, 77133334, 77199999}, '{A5, 77200000, 77495833}, '{PAUSE, 77495834, 77499999}, '{G5, 77500000, 77895833}, '{PAUSE, 77895834, 77899999}, '{E5, 77900000, 78333333}, '{PAUSE, 78333334, 78399999}, '{C5, 78400000, 78733333}, '{PAUSE, 78733334, 78799999}, '{D_s5, 78800000, 79133333}, '{PAUSE, 79133334, 79199999}, '{G5, 79200000, 79533333}, '{PAUSE, 79533334, 79599999}, '{A5, 79600000, 79933333}, '{PAUSE, 79933334, 79999999}, '{A_s5, 80000000, 80295833}, '{PAUSE, 80295834, 80299999}, '{A5, 80300000, 80695833}, '{PAUSE, 80695834, 80699999}, '{G5, 80700000, 81500000}, '{PAUSE, 81500001, 81599999}, '{G5, 81600000, 81933333}, '{PAUSE, 81933334, 81999999}, '{A5, 82000000, 82333333}, 
'{PAUSE, 82333334, 82399999}, '{F_s5, 82400000, 82733333}, '{PAUSE, 82733334, 82799999}, '{G5, 82800000, 83095833}, '{PAUSE, 83095834, 83099999}, 
'{E5, 83100000, 83495833}, '{PAUSE, 83495834, 83499999}, '{F_s5, 83500000, 83895833}, '{PAUSE, 83895834, 83899999}, '{E5, 83900000, 84295833}, '{PAUSE, 84295834, 84299999}, '{D_s5, 84300000, 84733333}, '{PAUSE, 84733334, 84799999}, '{G5, 84800000, 85133333}, '{PAUSE, 85133334, 85199999}, '{A5, 85200000, 85533333}, '{PAUSE, 85533334, 85599999}, '{F_s5, 85600000, 85933333}, '{PAUSE, 85933334, 85999999}, '{G5, 86000000, 86295833}, '{PAUSE, 86295834, 86299999}, '{E5, 86300000, 86695833}, '{PAUSE, 86695834, 86699999}, '{F_s5, 86700000, 87095833}, '{PAUSE, 87095834, 87099999}, '{D_s5, 87100000, 87533333}, '{PAUSE, 87533334, 87999999}, '{D5, 88000000, 88333333}, '{PAUSE, 88333334, 88399999}, '{E5, 88400000, 88733333}, '{PAUSE, 
88733334, 88799999}, '{G5, 88800000, 89133333}, '{PAUSE, 89133334, 89199999}, '{D6, 89200000, 89533333}, '{PAUSE, 89533334, 89599999}, '{C6, 89600000, 91100000}, '{PAUSE, 91100001, 91199999}, '{B5, 91200000, 91533333}, '{PAUSE, 91533334, 91599999}, '{A5, 91600000, 91933333}, '{PAUSE, 91933334, 91999999}, '{G5, 92000000, 92333333}, '{PAUSE, 92333334, 92399999}, '{E5, 92400000, 92733333}, '{PAUSE, 92733334, 92799999}, '{D_s5, 92800000, 
93133333}, '{PAUSE, 93133334, 93199999}, '{A5, 93200000, 93900000}, '{PAUSE, 93900001, 93999999}, '{B5, 94000000, 94333333}, '{PAUSE, 94333334, 94399999}, '{A5, 94400000, 94695833}, '{PAUSE, 94695834, 94699999}, '{G5, 94700000, 97500000}, '{PAUSE, 97500001, 100799999}, '{B5, 100800000, 101133333}, '{PAUSE, 101133334, 101199999}, '{A5, 101200000, 101533333}, '{PAUSE, 101533334, 101599999}, '{G5, 101600000, 101933333}, '{PAUSE, 101933334, 101999999}, '{F_s5, 102000000, 102295833}, '{PAUSE, 102295834, 102299999}, '{G5, 102300000, 102695833}, '{PAUSE, 102695834, 102699999}, '{F_s5, 102700000, 103095833}, '{PAUSE, 103095834, 103099999}, '{E5, 103100000, 103195833}, '{PAUSE, 103195834, 103499999}, '{D5, 103500000, 103933333}, 
'{PAUSE, 103933334, 103999999}, '{A5, 104000000, 104333333}, '{PAUSE, 104333334, 104399999}, '{G5, 104400000, 104733333}, '{PAUSE, 104733334, 104799999}, '{G5, 104800000, 105133333}, '{PAUSE, 105133334, 105199999}, '{F_s5, 105200000, 105495833}, '{PAUSE, 105495834, 105499999}, '{G5, 105500000, 105895833}, '{PAUSE, 105895834, 105899999}, '{F_s5, 105900000, 106295833}, '{PAUSE, 106295834, 106299999}, '{E5, 106300000, 107100000}, '{PAUSE, 107100001, 107599999}, '{B5, 107600000, 107895833}, '{PAUSE, 107895834, 107899999}, '{A5, 107900000, 107995833}, '{PAUSE, 107995834, 107999999}, '{A5, 108000000, 108295833}, '{PAUSE, 108295834, 108299999}, '{A5, 108300000, 108695833}, '{PAUSE, 108695834, 108699999}, '{B5, 108700000, 109095833}, '{PAUSE, 109095834, 109099999}, '{E6, 109100000, 109495833}, '{PAUSE, 109495834, 109499999}, '{A5, 109500000, 109895833}, '{PAUSE, 109895834, 109899999}, '{G5, 109900000, 110333333}, '{PAUSE, 110333334, 110799999}, '{B5, 110800000, 111095833}, '{PAUSE, 111095834, 111099999}, '{A5, 111100000, 111195833}, '{PAUSE, 111195834, 111199999}, '{B5, 111200000, 111495833}, '{PAUSE, 111495834, 111499999}, '{A5, 111500000, 111895833}, '{PAUSE, 111895834, 111899999}, '{B5, 111900000, 112295833}, '{PAUSE, 112295834, 112299999}, '{A5, 112300000, 112695833}, '{PAUSE, 112695834, 112699999}, '{G5, 112700000, 113500000}, '{PAUSE, 113500001, 113599999}, '{A5, 113600000, 113933333}, '{PAUSE, 113933334, 113999999}, '{G5, 114000000, 114295833}, '{PAUSE, 114295834, 114299999}, '{G5, 114300000, 114695833}, '{PAUSE, 114695834, 114699999}, '{F_s5, 114700000, 115095833}, '{PAUSE, 115095834, 115099999}, '{G5, 115100000, 115495833}, '{PAUSE, 115495834, 115499999}, '{F_s5, 115500000, 115895833}, '{PAUSE, 115895834, 115899999}, '{E5, 115900000, 116295833}, '{PAUSE, 116295834, 116299999}, '{D5, 116300000, 116733333}, '{PAUSE, 116733334, 116799999}, '{G4, 116800000, 117133333}, '{PAUSE, 117133334, 117199999}, '{B4, 117200000, 117495833}, '{PAUSE, 117495834, 117499999}, '{D5, 117500000, 117895833}, '{PAUSE, 117895834, 117899999}, '{F_s5, 117900000, 118295833}, '{PAUSE, 118295834, 118299999}, '{G5, 118300000, 118695833}, '{PAUSE, 118695834, 118699999}, '{F_s5, 118700000, 119095833}, '{PAUSE, 119095834, 119099999}, '{E5, 119100000, 119900000}, '{PAUSE, 119900001, 120399999}, '{B5, 120400000, 120695833}, '{PAUSE, 120695834, 120699999}, '{A5, 120700000, 120795833}, '{PAUSE, 120795834, 120799999}, '{B5, 120800000, 121095833}, '{PAUSE, 121095834, 121099999}, '{A5, 121100000, 121495833}, '{PAUSE, 121495834, 121499999}, '{B5, 121500000, 121895833}, '{PAUSE, 121895834, 121899999}, '{A5, 121900000, 122295833}, '{PAUSE, 122295834, 122299999}, '{G5, 122300000, 122695833}, '{PAUSE, 122695834, 122699999}, '{E5, 122700000, 123133333}, '{PAUSE, 123133334, 123199999}, '{C5, 123200000, 123533333}, '{PAUSE, 123533334, 123599999}, '{D_s5, 123600000, 123933333}, '{PAUSE, 123933334, 123999999}, '{G5, 124000000, 124333333}, '{PAUSE, 124333334, 124399999}, '{A5, 124400000, 124733333}, '{PAUSE, 124733334, 124799999}, '{A_s5, 124800000, 125095833}, 
'{PAUSE, 125095834, 125099999}, '{A5, 125100000, 125495833}, '{PAUSE, 125495834, 125499999}, '{G5, 125500000, 126295833}, '{PAUSE, 126295834, 126299999}, '{G5, 126300000, 126395833}, '{PAUSE, 126395834, 126399999}, '{G5, 126400000, 126733333}, '{PAUSE, 126733334, 126799999}, '{A5, 126800000, 127133333}, '{PAUSE, 127133334, 127199999}, '{F_s5, 127200000, 127533333}, '{PAUSE, 127533334, 127599999}, '{G5, 127600000, 127933333}, '{PAUSE, 
127933334, 127999999}, '{E5, 128000000, 128295833}, '{PAUSE, 128295834, 128299999}, '{F_s5, 128300000, 128695833}, '{PAUSE, 128695834, 128699999}, '{E5, 128700000, 129095833}, '{PAUSE, 129095834, 129099999}, '{D_s5, 129100000, 129533333}, '{PAUSE, 129533334, 129599999}, '{B5, 129600000, 129933333}, '{PAUSE, 129933334, 129999999}, '{A5, 130000000, 130333333}, '{PAUSE, 130333334, 130399999}, '{A5, 130400000, 130733333}, '{PAUSE, 130733334, 130799999}, '{G5, 130800000, 131133333}, '{PAUSE, 131133334, 131199999}, '{G5, 131200000, 131495833}, '{PAUSE, 131495834, 131499999}, '{A5, 131500000, 131895833}, '{PAUSE, 131895834, 131899999}, '{D_s5, 131900000, 132695833}, '{PAUSE, 132695834, 132699999}, '{D5, 132700000, 132795833}, '{PAUSE, 132795834, 132799999}, '{D5, 132800000, 133133333}, '{PAUSE, 133133334, 133199999}, '{E5, 133200000, 133533333}, '{PAUSE, 133533334, 133599999}, '{G5, 133600000, 133933333}, '{PAUSE, 133933334, 133999999}, '{D6, 134000000, 134333333}, '{PAUSE, 134333334, 134399999}, '{C6, 134400000, 
135100000}, '{PAUSE, 135100001, 135599999}, '{C6, 135600000, 135895833}, '{PAUSE, 135895834, 135899999}, '{D6, 135900000, 135995833}, '{PAUSE, 135995834, 135999999}, '{B5, 136000000, 136333333}, '{PAUSE, 136333334, 136399999}, '{A5, 136400000, 136733333}, '{PAUSE, 136733334, 136799999}, '{G5, 136800000, 137133333}, '{PAUSE, 137133334, 137199999}, '{E5, 137200000, 137533333}, '{PAUSE, 137533334, 137599999}, '{D_s5, 137600000, 137933333}, '{PAUSE, 137933334, 137999999}, '{A5, 138000000, 138700000}, '{PAUSE, 138700001, 138799999}, '{B5, 138800000, 139133333}, '{PAUSE, 139133334, 139199999}, '{G5, 139200000, 141900000}, '{PAUSE, 141900001, 146399999}, '{B5, 146400000, 146733333}, '{PAUSE, 146733334, 146799999}, '{B5, 146800000, 147095833}, '{PAUSE, 147095834, 147099999}, '{C6, 147100000, 147495833}, '{PAUSE, 147495834, 147499999}, '{B5, 147500000, 147895833}, '{PAUSE, 147895834, 147899999}, '{A5, 147900000, 148295833}, '{PAUSE, 148295834, 148299999}, '{G5, 148300000, 148695833}, '{PAUSE, 148695834, 148699999}, 
'{F_s5, 148700000, 148795833}, '{PAUSE, 148795834, 148799999}, '{E5, 148800000, 149133333}, '{PAUSE, 149133334, 149199999}, '{F_s5, 149200000, 149533333}, '{PAUSE, 149533334, 149599999}, '{G5, 149600000, 149933333}, '{PAUSE, 149933334, 149999999}, '{A5, 150000000, 150295833}, '{PAUSE, 150295834, 150299999}, '{G5, 150300000, 151100000}, '{PAUSE, 151100001, 152799999}, '{B5, 152800000, 153133333}, '{PAUSE, 153133334, 153199999}, '{B5, 153200000, 153495833}, '{PAUSE, 153495834, 153499999}, '{E6, 153500000, 153895833}, '{PAUSE, 153895834, 153899999}, '{D6, 153900000, 154295833}, '{PAUSE, 154295834, 154299999}, '{B5, 154300000, 154695833}, '{PAUSE, 154695834, 154699999}, '{A5, 154700000, 155133333}, '{PAUSE, 155133334, 155199999}, '{G5, 155200000, 155533333}, '{PAUSE, 155533334, 155599999}, '{A5, 155600000, 155933333}, '{PAUSE, 155933334, 155999999}, '{B5, 156000000, 156333333}, '{PAUSE, 156333334, 156399999}, '{A5, 156400000, 156695833}, '{PAUSE, 156695834, 156699999}, '{G5, 156700000, 157500000}, '{PAUSE, 157500001, 159099999}, '{G5, 159100000, 159195833}, '{PAUSE, 159195834, 159199999}, '{A5, 159200000, 159495833}, '{PAUSE, 159495834, 159499999}, '{A5, 159500000, 159895833}, '{PAUSE, 159895834, 159899999}, '{A5, 159900000, 160295833}, '{PAUSE, 160295834, 160299999}, '{A5, 160300000, 160695833}, 
'{PAUSE, 160695834, 160699999}, '{A5, 160700000, 161095833}, '{PAUSE, 161095834, 161099999}, '{G5, 161100000, 161933333}, '{PAUSE, 161933334, 162299999}, '{A5, 162300000, 162395833}, '{PAUSE, 162395834, 162399999}, '{B5, 162400000, 162695833}, '{PAUSE, 162695834, 162699999}, '{B5, 162700000, 163095833}, '{PAUSE, 163095834, 163099999}, '{E6, 163100000, 163495833}, '{PAUSE, 163495834, 163499999}, '{D6, 163500000, 163895833}, '{PAUSE, 163895834, 163899999}, '{B5, 163900000, 164295833}, '{PAUSE, 164295834, 164299999}, '{A5, 164300000, 164733333}, '{PAUSE, 164733334, 164799999}, '{B5, 164800000, 165095833}, '{PAUSE, 165095834, 165099999}, '{B5, 165100000, 165195833}, '{PAUSE, 165195834, 165199999}, '{B5, 165200000, 165495833}, '{PAUSE, 165495834, 165499999}, '{B5, 165500000, 165595833}, '{PAUSE, 165595834, 165599999}, '{B5, 165600000, 165933333}, '{PAUSE, 165933334, 165999999}, '{B5, 166000000, 166295833}, '{PAUSE, 166295834, 166299999}, '{B5, 166300000, 166395833}, '{PAUSE, 166395834, 166399999}, '{B5, 166400000, 166695833}, '{PAUSE, 166695834, 166699999}, '{B5, 166700000, 166795833}, '{PAUSE, 166795834, 166799999}, '{B5, 166800000, 167095833}, '{PAUSE, 
167095834, 167099999}, '{B5, 167100000, 167195833}, '{PAUSE, 167195834, 167199999}, '{B5, 167200000, 167533333}, '{PAUSE, 167533334, 167599999}, '{B5, 167600000, 167895833}, '{PAUSE, 167895834, 167899999}, '{B5, 167900000, 167995833}, '{PAUSE, 167995834, 167999999}, '{E6, 168000000, 168333333}, '{PAUSE, 168333334, 168399999}, '{D6, 168400000, 168733333}, '{PAUSE, 168733334, 168799999}, '{D6, 168800000, 169095833}, '{PAUSE, 169095834, 
169099999}, '{B5, 169100000, 169195833}, '{PAUSE, 169195834, 169199999}, '{D6, 169200000, 169495833}, '{PAUSE, 169495834, 169499999}, '{D6, 169500000, 169895833}, '{PAUSE, 169895834, 169899999}, '{B5, 169900000, 170333333}, '{PAUSE, 170333334, 171199999}, '{A5, 171200000, 171533333}, '{PAUSE, 171533334, 171599999}, '{G5, 171600000, 171933333}, '{PAUSE, 171933334, 171999999}, '{G5, 172000000, 172333333}, '{PAUSE, 172333334, 172399999}, '{F_s5, 172400000, 172695833}, '{PAUSE, 172695834, 172699999}, '{G5, 172700000, 173095833}, '{PAUSE, 173095834, 173099999}, '{F_s5, 173100000, 173495833}, '{PAUSE, 173495834, 173499999}, '{E5, 173500000, 173895833}, '{PAUSE, 173895834, 173899999}, '{D5, 173900000, 174333333}, '{PAUSE, 174333334, 174399999}, '{A5, 174400000, 174733333}, '{PAUSE, 174733334, 174799999}, '{G5, 174800000, 175133333}, '{PAUSE, 175133334, 175199999}, '{G5, 
175200000, 175533333}, '{PAUSE, 175533334, 175599999}, '{F_s5, 175600000, 175895833}, '{PAUSE, 175895834, 175899999}, '{G5, 175900000, 176295833}, '{PAUSE, 176295834, 176299999}, '{F_s5, 176300000, 176695833}, '{PAUSE, 176695834, 176699999}, '{E5, 176700000, 177500000}, '{PAUSE, 177500001, 177999999}, '{B5, 178000000, 178295833}, '{PAUSE, 178295834, 178299999}, '{A5, 178300000, 178395833}, '{PAUSE, 178395834, 178399999}, '{B5, 178400000, 178733333}, '{PAUSE, 178733334, 178799999}, '{A5, 178800000, 179095833}, '{PAUSE, 179095834, 179099999}, '{B5, 179100000, 179495833}, '{PAUSE, 179495834, 179499999}, '{E6, 179500000, 179895833}, '{PAUSE, 179895834, 179899999}, '{A5, 179900000, 180295833}, '{PAUSE, 180295834, 180299999}, 
'{G5, 180300000, 180733333}, '{PAUSE, 180733334, 180799999}, '{B5, 180800000, 181133333}, '{PAUSE, 181133334, 181199999}, '{A5, 181200000, 181495833}, '{PAUSE, 181495834, 181499999}, '{B5, 181500000, 181895833}, '{PAUSE, 181895834, 181899999}, '{A5, 181900000, 182295833}, '{PAUSE, 182295834, 182299999}, '{B5, 182300000, 182695833}, '{PAUSE, 182695834, 182699999}, '{A5, 182700000, 183095833}, '{PAUSE, 183095834, 183099999}, '{G5, 183100000, 183900000}, '{PAUSE, 183900001, 183999999}, '{G5, 184000000, 184333333}, '{PAUSE, 184333334, 184399999}, '{A5, 184400000, 184733333}, '{PAUSE, 184733334, 184799999}, '{F_s5, 184800000, 185133333}, '{PAUSE, 185133334, 185199999}, '{G5, 185200000, 185495833}, '{PAUSE, 185495834, 185499999}, '{E5, 185500000, 185895833}, '{PAUSE, 185895834, 185899999}, '{F_s5, 185900000, 186295833}, '{PAUSE, 186295834, 186299999}, '{E5, 186300000, 186695833}, '{PAUSE, 186695834, 186699999}, '{D_s5, 186700000, 187133333}, '{PAUSE, 187133334, 187199999}, '{G5, 187200000, 187533333}, '{PAUSE, 187533334, 187599999}, '{A5, 187600000, 187933333}, '{PAUSE, 187933334, 187999999}, '{F_s5, 188000000, 188333333}, '{PAUSE, 188333334, 188399999}, '{G5, 188400000, 188695833}, '{PAUSE, 188695834, 188699999}, '{E5, 188700000, 189095833}, '{PAUSE, 189095834, 189099999}, '{F_s5, 189100000, 189495833}, '{PAUSE, 189495834, 189499999}, '{D_s5, 189500000, 190300000}, '{PAUSE, 190300001, 190399999}, '{D5, 190400000, 190733333}, '{PAUSE, 190733334, 190799999}, '{E5, 190800000, 191133333}, '{PAUSE, 191133334, 191199999}, '{G5, 191200000, 191533333}, '{PAUSE, 191533334, 191599999}, '{D6, 191600000, 191933333}, '{PAUSE, 191933334, 191999999}, '{C6, 192000000, 193500000}, '{PAUSE, 193500001, 193599999}, '{B5, 193600000, 193933333}, '{PAUSE, 193933334, 193999999}, '{A5, 194000000, 194333333}, '{PAUSE, 194333334, 194399999}, '{G5, 194400000, 194733333}, '{PAUSE, 194733334, 194799999}, '{E5, 194800000, 195133333}, '{PAUSE, 195133334, 195199999}, '{D_s5, 195200000, 195533333}, '{PAUSE, 195533334, 195599999}, '{A5, 195600000, 
197500000}, '{PAUSE, 197500001, 197599999}, '{B5, 197600000, 198733333}, '{PAUSE, 198733334, 199999999}, '{G6, 200000000, 206300000}, '{PAUSE, 200000001, 202000001}};




module PIEZO_BGMUSIC (
    clk,
    dipswitch_two,
    music_idx,

    piezo
);


    initial begin
        cnt_piezo <= 0;
        cnt_piezo_two <= 0;
        cnt_piezo_three <= 0;

        piezo_bunzu <= 0;

        note_idx = 0;
        note_idx_two = 0;
        note_idx_three = 0;

        cur_tone = 3822;
        cur_start <= 0;
        cur_last <= 2147483647;
    end

    input wire clk;
    input wire dipswitch_two;
    input wire music_idx;

    output reg piezo;

    int note_idx, note_idx_two, note_idx_three;
    int cur_tone, cur_start, cur_last;
    int cnt_piezo, cnt_piezo_two, cnt_piezo_three;
    int piezo_bunzu;

    always @(posedge clk) begin
        if (dipswitch_two == 1'b1) begin
            if (music_idx == 2'b00) begin

                if (cur_start <= cnt_piezo && cnt_piezo <= cur_last) begin
                    if (cur_tone == PAUSE) begin
                    end

                    else if (cur_tone == ENDL) begin
                        note_idx = 0;
                        cnt_piezo = -1;
                        // Reset to the first note of the tune
                        cur_tone = ballgame[0].tone;
                        cur_start = ballgame[0].sstart;
                        cur_last = ballgame[0].llast;
                    end

                    else if (piezo_bunzu >= cur_tone/2) begin
                        piezo = !piezo;
                        piezo_bunzu = 0;
                    end

                    else begin
                        piezo_bunzu = piezo_bunzu + 1;
                    end
                end

                else begin
                    note_idx <= (note_idx + 1);
                    cur_tone <= ballgame[note_idx].tone;
                    cur_start <= ballgame[note_idx].sstart;
                    cur_last <= ballgame[note_idx].llast;
                end
                
                cnt_piezo = cnt_piezo + 1;
            end

            else if (music_idx == 1) begin
                if (cur_start <= cnt_piezo_two && cnt_piezo_two <= cur_last) begin
                    if (cur_tone == PAUSE) begin
                    end
                    
                    else if (piezo_bunzu >= cur_tone/2) begin
                        piezo = !piezo;
                        piezo_bunzu = 0;
                    end

                    else begin
                        piezo_bunzu = piezo_bunzu + 1;
                    end
                end

                else begin
                    note_idx_two <= (note_idx_two + 1);
                    cur_tone <= dearX[note_idx_two].tone;
                    cur_start <= dearX[note_idx_two].sstart;
                    cur_last <= dearX[note_idx_two].llast;
                end

                cnt_piezo_two = cnt_piezo_two + 1;

            end

            else if (music_idx == 2) begin
                if (cur_start <= cnt_piezo_three && cnt_piezo_three <= cur_last) begin

                    if (cur_tone == PAUSE) begin
                    end

                    else if (piezo_bunzu >= cur_tone/2) begin
                        piezo = !piezo;
                        piezo_bunzu = 0;
                    end

                    else begin
                        piezo_bunzu = piezo_bunzu + 1;
                    end
                end

                else begin
                    note_idx_three <= (note_idx_three + 1);
                    cur_tone <= narco[note_idx_three].tone;
                    cur_start <= narco[note_idx_three].sstart;
                    cur_last <= narco[note_idx_three].llast;
                end

                cnt_piezo_three = cnt_piezo_three + 1;
            end
        end

        else begin // dipswitch_two == 1'b0
            note_idx = 0;
            note_idx_two = 0;
            note_idx_three = 0;
            cur_tone = ballgame[0].tone;
            cur_start = ballgame[0].sstart;
            cur_last = ballgame[0].llast;
            cnt_piezo_two = 0;
            cnt_piezo = 0;
        end
    end

endmodule
